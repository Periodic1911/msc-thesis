module alu(
  input logic [3:0] ALUControlE,
  input logic [31:0] Op1E, Op2E,

  output logic [31:0] ALUResultE,
  output logic [3:0] ALUFlags, // ARM only
  output logic ZeroE // RISC-V only
);

logic [31:0] addResult;

add_sub as(.a(Op1E), .b(Op2E), .q(addResult), .add(~ALUControlE[0]), .cOut(carry),
  .overflow(overflow) // ARM only
  );

logic [31:0] shiftResult;

barrel_shift bs(Op1E, Op2E[4:0], shiftOp, shiftResult);

always_comb
  case(ALUControlE)
    4'b0000: ALUResultE = addResult; // add
    4'b0001: ALUResultE = addResult; // sub
    4'b0010: ALUResultE = Op1E & Op2E; // and
    4'b0011: ALUResultE = Op1E | Op2E; // or
    4'b0100: ALUResultE = Op1E ^ Op2E; // xor
    // RISC-V only
    4'b0101: ALUResultE = (Op1E < Op2E) ? 32'b1 : 32'b0; // slt TODO: reuse add_sub carry chain?
    default: ALUResultE = 32'hxxxxxxxx; /// ???
  endcase

assign ZeroE = (ALUResultE == 0); // RISC-V only

logic neg, zero, carry, overflow; // ARM only
assign ALUFlags = {neg, zero, carry, overflow}; // ARM only

always_comb begin : ARM_Flags // ARM only
  zero = (ALUResultE == 0);
  neg = ALUResultE[31];
end

endmodule

/* Combined adder-subtractor with one carry chain */
module add_sub(
  input logic [31:0] a, b,
  input logic add,
  output logic [31:0] q,
  output logic cOut,
  output logic overflow // ARM only
);

logic [31:0] b_inv;
assign b_inv = add ? b : ~b;
logic carry_in = ~add;
logic carry_out;

assign {carry_out, q} = a + b_inv + {31'b0, carry_in};
xor(cOut, carry_out, carry_in);
assign overflow = (~q[31] & a[31] & b_inv[31]) |
                  ( q[31] &~a[31] &~b_inv[31]);

endmodule

/* Barrel shifter with support for
* - 00 logical left shift
* - 10/01 arithmetic/logical right shift
* - 11 rotate right
*/
module barrel_shift(
  input logic [31:0] a,
  input logic [4:0] shift,
  input logic [1:0] op,
  output logic [31:0] q
);

logic signExt;
assign signExt = (op == 2'b10) ? a[31] : 1'b0;
logic rot = (op == 2'b11);

logic [31:0] arshift_stage [4:0];
mux2 #(32) barshift16 (a, {{16{signExt}}, a[31:16]}, shift[4], arshift_stage[4]);
mux2 #(32) barshift8 (arshift_stage[4], {{8{signExt}}, arshift_stage[4][31:8]}, shift[3], arshift_stage[3]);
mux2 #(32) barshift4 (arshift_stage[3], {{4{signExt}}, arshift_stage[3][31:4]}, shift[2], arshift_stage[2]);
mux2 #(32) barshift2 (arshift_stage[2], {{2{signExt}}, arshift_stage[2][31:2]}, shift[1], arshift_stage[1]);
mux2 #(32) barshift1 (arshift_stage[1], {signExt, arshift_stage[1][31:1]}, shift[0], arshift_stage[0]);

logic [31:0] ror_stage [4:0];
mux2 #(32) bror16 (a, {a[15:0], a[31:16]}, shift[4], ror_stage[4]);
mux2 #(32) bror8 (ror_stage[4], {ror_stage[4][7:0], ror_stage[4][31:8]}, shift[3], ror_stage[3]);
mux2 #(32) bror4 (ror_stage[3], {ror_stage[3][3:0], ror_stage[3][31:4]}, shift[2], ror_stage[2]);
mux2 #(32) bror2 (ror_stage[2], {ror_stage[2][1:0], ror_stage[2][31:2]}, shift[1], ror_stage[1]);
mux2 #(32) bror1 (ror_stage[1], {ror_stage[1][0], ror_stage[1][31:1]}, shift[0], ror_stage[0]);

logic [31:0] lshift_stage [4:0];
mux2 #(32) blshift16 (a, {a[15:0], 16'b0}, shift[4], lshift_stage[4]);
mux2 #(32) blshift8 (lshift_stage[4], {lshift_stage[4][23:0], 8'b0}, shift[3], lshift_stage[3]);
mux2 #(32) blshift4 (lshift_stage[3], {lshift_stage[3][27:0], 4'b0}, shift[2], lshift_stage[2]);
mux2 #(32) blshift2 (lshift_stage[2], {lshift_stage[2][29:0], 2'b0}, shift[1], lshift_stage[1]);
mux2 #(32) blshift1 (lshift_stage[1], {lshift_stage[1][30:0], 1'b0}, shift[0], lshift_stage[0]);

always_comb
  case(op)
    2'b00: q = lshift_stage[0];
    2'b01: q = arshift_stage[0];
    2'b10: q = arshift_stage[0];
    2'b11: q = ror_stage[0];
  endcase

endmodule
